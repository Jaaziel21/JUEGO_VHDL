-- Contador de pixeles (525) en el plano vertical para un esquema de 640x480 pixeles
-- Leyberth Jaaziel Castillo Guerra	A01749505
-- Maximiliano De La Cruz Lima	A01798048
-- TE2002B

-- Librerías
library ieee;
use ieee.std_logic_1164.all;

-- Definición de la entidad
entity contador500 is
	
	port ( CLK, RST, START : in std_logic;						-- Entradas
			 CNT : out std_logic_vector (9 downto 0);	-- Salidas
			 OVout : out std_logic);
			 
end entity;

architecture RTL of contador500 is
	
	-- Definición de los componentes
		
			-- Definición del uso de componente SUMA_10BITS
			
			component mas_uno_10bits is
				
				port ( A		: in 	std_logic_vector (9 downto 0);	-- Entradas
						 Z		: out std_logic_vector (9 downto 0);	-- Salidas
						 Cout	: out std_logic );
				
			end component mas_uno_10bits;
	
	-- Cables de interconexión
		
	signal D, Q 		: std_logic_vector (9 downto 0);
	signal O	: std_logic;

	-- Descripción del circuito
	
	begin
	
		SUMA10 : mas_uno_10bits port map ( Q, D, O );
			
					FFD : process (CLK, RST)
			
				begin
				
					if (RST = '0') then
						Q <= "0000000000";
						OVout <= '0';
					elsif (CLK'EVENT and CLK = '1') then
						if (START = '1') then
							Q <= D;
						end if;
						if (Q = "1000001100") then
							Q <= "0000000000";
							OVout <= '1';
						else
							OVout <= '0';
						end if;
					end if;
					
			end process FFD;	
			
			CNT <= Q;	
		
	
end architecture;